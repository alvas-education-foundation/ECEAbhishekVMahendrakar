<circuit>
<CurrentPage>0</CurrentPage>
<page 0>
<PageViewport>-7.75495,4.08436,96.795,-48.5656</PageViewport>
<gate>
<ID>2</ID>
<type>AA_MUX_2x1</type>
<position>14,-20.5</position>
<input>
<ID>IN_0</ID>9 </input>
<input>
<ID>IN_1</ID>8 </input>
<output>
<ID>OUT</ID>10 </output>
<input>
<ID>SEL_0</ID>2 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>4</ID>
<type>AA_TOGGLE</type>
<position>8,-5</position>
<output>
<ID>OUT_0</ID>2 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>6</ID>
<type>AA_TOGGLE</type>
<position>23.5,-5</position>
<output>
<ID>OUT_0</ID>4 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>8</ID>
<type>AA_TOGGLE</type>
<position>37.5,-5</position>
<output>
<ID>OUT_0</ID>5 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>10</ID>
<type>AA_TOGGLE</type>
<position>60.5,-5.5</position>
<output>
<ID>OUT_0</ID>22 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>12</ID>
<type>GA_LED</type>
<position>74,-30</position>
<input>
<ID>N_in0</ID>29 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>14</ID>
<type>AA_MUX_2x1</type>
<position>27.5,-14</position>
<input>
<ID>IN_0</ID>7 </input>
<input>
<ID>IN_1</ID>12 </input>
<output>
<ID>OUT</ID>8 </output>
<input>
<ID>SEL_0</ID>4 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>16</ID>
<type>AA_MUX_2x1</type>
<position>32,-23.5</position>
<input>
<ID>IN_0</ID>5 </input>
<input>
<ID>IN_1</ID>11 </input>
<output>
<ID>OUT</ID>19 </output>
<input>
<ID>SEL_0</ID>10 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>18</ID>
<type>AA_MUX_2x1</type>
<position>32.5,-33.5</position>
<input>
<ID>IN_0</ID>5 </input>
<input>
<ID>IN_1</ID>6 </input>
<output>
<ID>OUT</ID>13 </output>
<input>
<ID>SEL_0</ID>2 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>20</ID>
<type>AA_MUX_2x1</type>
<position>44,-14.5</position>
<input>
<ID>IN_0</ID>23 </input>
<input>
<ID>IN_1</ID>22 </input>
<output>
<ID>OUT</ID>24 </output>
<input>
<ID>SEL_0</ID>4 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>22</ID>
<type>AA_MUX_2x1</type>
<position>47.5,-21</position>
<input>
<ID>IN_0</ID>26 </input>
<input>
<ID>IN_1</ID>25 </input>
<output>
<ID>OUT</ID>27 </output>
<input>
<ID>SEL_0</ID>24 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>24</ID>
<type>AA_MUX_2x1</type>
<position>53.5,-26</position>
<input>
<ID>IN_0</ID>28 </input>
<input>
<ID>IN_1</ID>27 </input>
<output>
<ID>OUT</ID>18 </output>
<input>
<ID>SEL_0</ID>19 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>26</ID>
<type>AA_MUX_2x1</type>
<position>67.5,-30</position>
<input>
<ID>IN_0</ID>16 </input>
<input>
<ID>IN_1</ID>17 </input>
<output>
<ID>OUT</ID>29 </output>
<input>
<ID>SEL_0</ID>18 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>28</ID>
<type>AA_MUX_2x1</type>
<position>63.5,-37.5</position>
<input>
<ID>IN_0</ID>15 </input>
<input>
<ID>IN_1</ID>14 </input>
<output>
<ID>OUT</ID>16 </output>
<input>
<ID>SEL_0</ID>13 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>32</ID>
<type>EE_VDD</type>
<position>26,-34.5</position>
<output>
<ID>OUT_0</ID>6 </output>
<gparam>angle 180</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>34</ID>
<type>EE_VDD</type>
<position>23,-17.5</position>
<output>
<ID>OUT_0</ID>7 </output>
<gparam>angle 180</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>36</ID>
<type>FF_GND</type>
<position>10.5,-24</position>
<output>
<ID>OUT_0</ID>9 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>38</ID>
<type>EE_VDD</type>
<position>26,-25</position>
<output>
<ID>OUT_0</ID>11 </output>
<gparam>angle 180</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>40</ID>
<type>FF_GND</type>
<position>20.5,-16</position>
<output>
<ID>OUT_0</ID>12 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>42</ID>
<type>FF_GND</type>
<position>56,-39.5</position>
<output>
<ID>OUT_0</ID>14 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>44</ID>
<type>EE_VDD</type>
<position>59.5,-40.5</position>
<output>
<ID>OUT_0</ID>15 </output>
<gparam>angle 180</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>46</ID>
<type>EE_VDD</type>
<position>62,-30.5</position>
<output>
<ID>OUT_0</ID>17 </output>
<gparam>angle 180</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>52</ID>
<type>FF_GND</type>
<position>40.5,-18.5</position>
<output>
<ID>OUT_0</ID>23 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>54</ID>
<type>FF_GND</type>
<position>40,-22</position>
<output>
<ID>OUT_0</ID>25 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>56</ID>
<type>EE_VDD</type>
<position>43,-25.5</position>
<output>
<ID>OUT_0</ID>26 </output>
<gparam>angle 180</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>58</ID>
<type>FF_GND</type>
<position>49.5,-29.5</position>
<output>
<ID>OUT_0</ID>28 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>60</ID>
<type>AA_LABEL</type>
<position>8,-2.5</position>
<gparam>LABEL_TEXT A</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>62</ID>
<type>AA_LABEL</type>
<position>23.5,-2.5</position>
<gparam>LABEL_TEXT B</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>64</ID>
<type>AA_LABEL</type>
<position>37.5,-2.5</position>
<gparam>LABEL_TEXT C</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>66</ID>
<type>AA_LABEL</type>
<position>60.5,-3</position>
<gparam>LABEL_TEXT D</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>68</ID>
<type>AA_LABEL</type>
<position>45,1</position>
<gparam>LABEL_TEXT Implementing Y = ( A.B '+ C ) . ((B.D)') + ( (A+C)') only using 2:1 MUX</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>70</ID>
<type>AA_LABEL</type>
<position>76.5,-29.5</position>
<gparam>LABEL_TEXT Y</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>74</ID>
<type>AA_LABEL</type>
<position>76.5,-43</position>
<gparam>LABEL_TEXT Name: Abhishek Vasudev Mahendrakar</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>76</ID>
<type>AA_LABEL</type>
<position>68.5,-45</position>
<gparam>LABEL_TEXT USN: 4AL17EC003</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>78</ID>
<type>AA_LABEL</type>
<position>68,-47</position>
<gparam>LABEL_TEXT SEM/SEC: 6th-'A'</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<wire>
<ID>2</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>8,-31,8,-7</points>
<connection>
<GID>4</GID>
<name>OUT_0</name></connection>
<intersection>-31 5</intersection>
<intersection>-12 6</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>8,-31,32.5,-31</points>
<connection>
<GID>18</GID>
<name>SEL_0</name></connection>
<intersection>8 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>8,-12,14,-12</points>
<intersection>8 0</intersection>
<intersection>14 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>14,-18,14,-12</points>
<connection>
<GID>2</GID>
<name>SEL_0</name></connection>
<intersection>-12 6</intersection></vsegment></shape></wire>
<wire>
<ID>4</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>27.5,-11.5,27.5,-8.5</points>
<connection>
<GID>14</GID>
<name>SEL_0</name></connection>
<intersection>-8.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>23.5,-8.5,23.5,-7</points>
<connection>
<GID>6</GID>
<name>OUT_0</name></connection>
<intersection>-8.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>23.5,-8.5,44,-8.5</points>
<intersection>23.5 1</intersection>
<intersection>27.5 0</intersection>
<intersection>44 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>44,-12,44,-8.5</points>
<connection>
<GID>20</GID>
<name>SEL_0</name></connection>
<intersection>-8.5 2</intersection></vsegment></shape></wire>
<wire>
<ID>5</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>37.5,-26.5,37.5,-7</points>
<connection>
<GID>8</GID>
<name>OUT_0</name></connection>
<intersection>-26.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>28,-26.5,37.5,-26.5</points>
<intersection>28 2</intersection>
<intersection>37.5 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>28,-34.5,28,-24.5</points>
<intersection>-34.5 4</intersection>
<intersection>-26.5 1</intersection>
<intersection>-24.5 5</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>28,-34.5,30.5,-34.5</points>
<connection>
<GID>18</GID>
<name>IN_0</name></connection>
<intersection>28 2</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>28,-24.5,30,-24.5</points>
<connection>
<GID>16</GID>
<name>IN_0</name></connection>
<intersection>28 2</intersection></hsegment></shape></wire>
<wire>
<ID>6</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>26,-33.5,26,-32.5</points>
<connection>
<GID>32</GID>
<name>OUT_0</name></connection>
<intersection>-32.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>26,-32.5,30.5,-32.5</points>
<connection>
<GID>18</GID>
<name>IN_1</name></connection>
<intersection>26 0</intersection></hsegment></shape></wire>
<wire>
<ID>7</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>23,-16.5,23,-15</points>
<connection>
<GID>34</GID>
<name>OUT_0</name></connection>
<intersection>-15 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>23,-15,25.5,-15</points>
<connection>
<GID>14</GID>
<name>IN_0</name></connection>
<intersection>23 0</intersection></hsegment></shape></wire>
<wire>
<ID>8</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>12,-10.5,29.5,-10.5</points>
<intersection>12 3</intersection>
<intersection>29.5 4</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>12,-19.5,12,-10.5</points>
<connection>
<GID>2</GID>
<name>IN_1</name></connection>
<intersection>-10.5 1</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>29.5,-14,29.5,-10.5</points>
<connection>
<GID>14</GID>
<name>OUT</name></connection>
<intersection>-10.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>9</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>10.5,-23,10.5,-21.5</points>
<connection>
<GID>36</GID>
<name>OUT_0</name></connection>
<intersection>-21.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>10.5,-21.5,12,-21.5</points>
<connection>
<GID>2</GID>
<name>IN_0</name></connection>
<intersection>10.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>10</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>32,-21,32,-20.5</points>
<connection>
<GID>16</GID>
<name>SEL_0</name></connection>
<intersection>-20.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>16,-20.5,32,-20.5</points>
<connection>
<GID>2</GID>
<name>OUT</name></connection>
<intersection>32 0</intersection></hsegment></shape></wire>
<wire>
<ID>11</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>26,-22.5,30,-22.5</points>
<connection>
<GID>16</GID>
<name>IN_1</name></connection>
<intersection>26 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>26,-24,26,-22.5</points>
<connection>
<GID>38</GID>
<name>OUT_0</name></connection>
<intersection>-22.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>12</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>20.5,-15,20.5,-13</points>
<connection>
<GID>40</GID>
<name>OUT_0</name></connection>
<intersection>-13 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>20.5,-13,25.5,-13</points>
<connection>
<GID>14</GID>
<name>IN_1</name></connection>
<intersection>20.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>13</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>63.5,-35,63.5,-33.5</points>
<connection>
<GID>28</GID>
<name>SEL_0</name></connection>
<intersection>-33.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>34.5,-33.5,63.5,-33.5</points>
<connection>
<GID>18</GID>
<name>OUT</name></connection>
<intersection>63.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>14</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>56,-38.5,56,-36.5</points>
<connection>
<GID>42</GID>
<name>OUT_0</name></connection>
<intersection>-36.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>56,-36.5,61.5,-36.5</points>
<connection>
<GID>28</GID>
<name>IN_1</name></connection>
<intersection>56 0</intersection></hsegment></shape></wire>
<wire>
<ID>15</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>59.5,-38.5,61.5,-38.5</points>
<connection>
<GID>28</GID>
<name>IN_0</name></connection>
<intersection>59.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>59.5,-39.5,59.5,-38.5</points>
<connection>
<GID>44</GID>
<name>OUT_0</name></connection>
<intersection>-38.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>16</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>65.5,-37.5,65.5,-31</points>
<connection>
<GID>26</GID>
<name>IN_0</name></connection>
<connection>
<GID>28</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>17</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>62,-29.5,62,-29</points>
<connection>
<GID>46</GID>
<name>OUT_0</name></connection>
<intersection>-29 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>62,-29,65.5,-29</points>
<connection>
<GID>26</GID>
<name>IN_1</name></connection>
<intersection>62 0</intersection></hsegment></shape></wire>
<wire>
<ID>18</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>67.5,-27.5,67.5,-26</points>
<connection>
<GID>26</GID>
<name>SEL_0</name></connection>
<intersection>-26 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>55.5,-26,67.5,-26</points>
<connection>
<GID>24</GID>
<name>OUT</name></connection>
<intersection>67.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>19</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>34,-23.5,53.5,-23.5</points>
<connection>
<GID>16</GID>
<name>OUT</name></connection>
<intersection>53.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>53.5,-23.5,53.5,-23.5</points>
<connection>
<GID>24</GID>
<name>SEL_0</name></connection>
<intersection>-23.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>22</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>60.5,-11,60.5,-7.5</points>
<connection>
<GID>10</GID>
<name>OUT_0</name></connection>
<intersection>-11 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>42,-11,60.5,-11</points>
<intersection>42 2</intersection>
<intersection>60.5 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>42,-13.5,42,-11</points>
<connection>
<GID>20</GID>
<name>IN_1</name></connection>
<intersection>-11 1</intersection></vsegment></shape></wire>
<wire>
<ID>23</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>40.5,-17.5,40.5,-15.5</points>
<connection>
<GID>52</GID>
<name>OUT_0</name></connection>
<intersection>-15.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>40.5,-15.5,42,-15.5</points>
<connection>
<GID>20</GID>
<name>IN_0</name></connection>
<intersection>40.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>24</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>47.5,-18.5,47.5,-14.5</points>
<connection>
<GID>22</GID>
<name>SEL_0</name></connection>
<intersection>-14.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>46,-14.5,47.5,-14.5</points>
<connection>
<GID>20</GID>
<name>OUT</name></connection>
<intersection>47.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>25</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>40,-21,40,-20</points>
<connection>
<GID>54</GID>
<name>OUT_0</name></connection>
<intersection>-20 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>40,-20,45.5,-20</points>
<connection>
<GID>22</GID>
<name>IN_1</name></connection>
<intersection>40 0</intersection></hsegment></shape></wire>
<wire>
<ID>26</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>43,-24.5,43,-22</points>
<connection>
<GID>56</GID>
<name>OUT_0</name></connection>
<intersection>-22 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>43,-22,45.5,-22</points>
<connection>
<GID>22</GID>
<name>IN_0</name></connection>
<intersection>43 0</intersection></hsegment></shape></wire>
<wire>
<ID>27</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>50.5,-25,50.5,-21</points>
<intersection>-25 1</intersection>
<intersection>-21 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>50.5,-25,51.5,-25</points>
<connection>
<GID>24</GID>
<name>IN_1</name></connection>
<intersection>50.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>49.5,-21,50.5,-21</points>
<connection>
<GID>22</GID>
<name>OUT</name></connection>
<intersection>50.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>28</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>49.5,-28.5,49.5,-27</points>
<connection>
<GID>58</GID>
<name>OUT_0</name></connection>
<intersection>-27 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>49.5,-27,51.5,-27</points>
<connection>
<GID>24</GID>
<name>IN_0</name></connection>
<intersection>49.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>29</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>69.5,-30,73,-30</points>
<connection>
<GID>26</GID>
<name>OUT</name></connection>
<connection>
<GID>12</GID>
<name>N_in0</name></connection></hsegment></shape></wire></page 0>
<page 1>
<PageViewport>0,0,139.4,-70.2</PageViewport></page 1>
<page 2>
<PageViewport>0,0,139.4,-70.2</PageViewport></page 2>
<page 3>
<PageViewport>0,0,139.4,-70.2</PageViewport></page 3>
<page 4>
<PageViewport>0,0,139.4,-70.2</PageViewport></page 4>
<page 5>
<PageViewport>0,0,139.4,-70.2</PageViewport></page 5>
<page 6>
<PageViewport>0,0,139.4,-70.2</PageViewport></page 6>
<page 7>
<PageViewport>0,0,139.4,-70.2</PageViewport></page 7>
<page 8>
<PageViewport>0,0,139.4,-70.2</PageViewport></page 8>
<page 9>
<PageViewport>0,0,139.4,-70.2</PageViewport></page 9></circuit>